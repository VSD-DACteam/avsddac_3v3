magic
tech scmos
timestamp 1594222475
<< metal1 >>
rect 1851 1506 1880 1509
rect 215 1494 219 1500
rect 229 1494 236 1503
rect 1664 1499 1697 1503
rect 1875 1500 1880 1506
rect 1664 1461 1669 1499
rect 1956 1478 1958 1481
rect 1881 1473 1883 1477
rect 1878 1460 1880 1463
rect 2890 572 2895 576
<< m2contact >>
rect 1846 1506 1851 1510
rect 33 1500 40 1504
rect 210 1494 215 1500
rect 1122 1485 1127 1490
rect 2788 1485 2792 1490
rect 1664 1455 1669 1461
rect 1873 1460 1878 1465
rect 1224 572 1231 576
<< metal2 >>
rect 1837 1507 1846 1510
rect 40 1500 208 1503
rect 203 1494 210 1500
rect 215 1494 216 1500
rect 2788 1490 2792 1491
rect 1873 1465 1878 1466
rect 1878 1460 1880 1463
rect 1664 1453 1669 1455
rect 1231 573 1234 576
<< m3contact >>
rect 1832 1506 1837 1510
rect 1122 1490 1127 1495
rect 2788 1491 2792 1496
rect 1873 1466 1878 1471
rect 1664 1447 1669 1453
rect 1234 572 1239 576
<< metal3 >>
rect 1822 1507 1832 1510
rect 2788 1496 2792 1497
rect 1873 1471 1878 1472
rect 1664 1445 1669 1447
rect 1239 572 1242 576
<< m4contact >>
rect 1817 1506 1822 1510
rect 1122 1495 1127 1500
rect 2788 1497 2792 1502
rect 1873 1472 1878 1477
rect 1664 1439 1670 1445
rect 1242 572 1247 576
<< metal4 >>
rect 1807 1507 1817 1510
rect 1126 1500 1127 1503
rect 2499 1502 2791 1505
rect 1873 1477 1878 1478
rect 1664 575 1668 1439
rect 1247 572 1668 575
<< m5contact >>
rect 1802 1506 1807 1510
rect 1121 1500 1126 1505
rect 2494 1501 2499 1505
rect 1873 1478 1878 1485
<< metal5 >>
rect 1121 1507 1802 1510
rect 1121 1505 1127 1507
rect 1126 1500 1127 1505
rect 1872 1502 2494 1505
rect 1872 1486 1875 1502
rect 2499 1502 2501 1505
rect 1872 1485 1878 1486
rect 1872 1482 1873 1485
<< pseudo_rpoly >>
rect 1234 572 1239 576
rect 2890 572 2891 576
use resistor3  resistor3_0
timestamp 1594222023
transform -1 0 218 0 1 1487
box -15 6 2 14
use 9bitres  9bitres_0
timestamp 1594222023
transform 1 0 0 0 1 0
box 0 0 1663 1510
use vsdswitch  vsdswitch_0
timestamp 1594101072
transform 1 0 1874 0 1 1481
box 1 -21 83 22
use 9bitres  9bitres_1
timestamp 1594222023
transform 1 0 1666 0 1 0
box 0 0 1663 1510
<< labels >>
rlabel metal1 1881 1473 1881 1477 1 D9!
rlabel metal1 1958 1478 1958 1481 1 out_ten
rlabel metal1 2893 574 2893 574 1 gnd!
rlabel metal1 229 1503 236 1503 1 vref
<< end >>
