magic
tech scmos
timestamp 1594105324
<< metal1 >>
rect 102 133 106 157
rect 97 130 106 133
rect 105 108 106 111
rect 25 103 31 107
rect -73 82 -68 95
rect 95 90 106 93
rect 103 62 106 90
use vsdswitch  vsdswitch_0
timestamp 1594101072
transform 1 0 22 0 1 111
box 1 -21 83 22
use 2bitres  2bitres_0
timestamp 1594105324
transform 1 0 -76 0 1 110
box -15 -20 182 69
use 2bitres  2bitres_1
timestamp 1594105324
transform 1 0 -76 0 1 18
box -15 -20 182 69
<< labels >>
rlabel metal1 25 103 25 107 1 D2!
rlabel metal1 106 108 106 111 7 out_three
<< end >>
