magic
tech scmos
timestamp 1594209536
<< metal1 >>
rect 1125 1485 1126 1488
rect 1049 1480 1050 1484
rect 1223 572 1224 576
<< m2contact >>
rect 858 1504 863 1509
rect 1114 1506 1119 1510
rect 1044 1466 1048 1470
rect 1448 733 1453 737
rect 616 727 620 732
rect 384 566 390 571
<< metal2 >>
rect 840 1504 858 1509
rect 1119 1506 1120 1510
rect 1449 737 1452 740
rect 390 566 394 570
<< m3contact >>
rect 834 1504 840 1509
rect 1120 1506 1127 1510
rect 1039 1466 1044 1470
rect 1448 740 1453 745
rect 616 732 620 737
rect 394 566 400 570
<< metal3 >>
rect 1127 1506 1129 1510
rect 834 1503 839 1504
rect 814 1500 839 1503
rect 1035 1463 1039 1465
rect 616 737 619 761
rect 1449 745 1452 772
<< m4contact >>
rect 1129 1506 1135 1510
rect 805 1499 814 1503
rect 1035 1465 1039 1470
rect 1449 772 1454 776
rect 616 761 621 765
rect 400 566 406 570
<< metal4 >>
rect 1135 1507 1452 1510
rect 409 1500 805 1503
rect 409 569 412 1500
rect 1035 1462 1039 1465
rect 616 1459 1039 1462
rect 616 765 619 1459
rect 1449 776 1452 1507
rect 406 566 412 569
use 8bitres  8bitres_0
timestamp 1594209536
transform 1 0 0 0 1 754
box 0 -754 830 750
use vsdswitch  vsdswitch_0
timestamp 1594101072
transform 1 0 1042 0 1 1488
box 1 -21 83 22
use 8bitres  8bitres_1
timestamp 1594209536
transform 1 0 833 0 1 760
box 0 -754 830 750
<< labels >>
rlabel metal1 1126 1485 1126 1488 1 out_nine
rlabel metal1 1049 1480 1049 1484 1 D8!
rlabel metal1 1224 572 1224 576 1 res_out_9
<< end >>
